module spi(
    input wire clk,
    input wire slk,
    input wire pico,
    input wire cs,
    output wire[7:0] data,
    output wire data_ready
);

// TODO

endmodule