module seven_segment(input wire[3:0] binary,
                            output reg[7:0] out);
/**
 * 7 segment code converter
 */
endmodule
