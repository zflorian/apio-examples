module seven_segment_logic(input wire[3:0] x,
                            output wire A,
                            output wire B,
                            output wire C,
                            output wire D,
                            output wire E,
                            output wire F,
                            output wire G,
                            output wire DP);

// 1. Wahrheitstabelle aufstellen
// 2a. Schaltung aus Mintermen herleiten
// 2b. Schaltung aus Maxtermen herleiten                            

endmodule